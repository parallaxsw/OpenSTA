module square_bracket (
  \in[0].test ,
  \out[0].test 
);
  input \in[0].test ;
  wire \in[0].test ;

  output \out[0].test ;
  wire \out[0].test ;

  BUFx2_ASAP7_75t_R inst0 (
    .A( \in[0].test ),
    .Y( \out[0].test )
  );
endmodule